/**
 * Модуль: video_wb_master
 * Описание: Wishbone Master для видеоконтроллера.
 *            Читает данные из памяти по адресу, когда видеоконтроллер требует пиксель.
 *            Реализует простейший конечный автомат для управления шиной.
 *            Имеет высший приоритет при подключении к арбитру.
 *
 * Входы:
 *   clk          - Тактовая частота (должна быть синхронна с шиной и памятью)
 *   rst          - Сброс (активный уровень high)
 *   pixel_enable - Сигнал от генератора таймингов: '1' означает, что требуется загрузка нового пикселя.
 *   phys_addr    - 24-битный физический адрес для чтения, сформированный vid_addr_gen.
 *   wb_dat_i     - 8-битные данные, читаемые из шины Wishbone
 *   wb_ack_i     - Подтверждение операции от slave (памяти)
 *
 * Выходы:
 *   wb_cyc_o     - Сигнал начала цикла шины Wishbone
 *   wb_stb_o     - Строб данных (импульсный сигнал запроса)
 *   wb_adr_o     - 24-битный адрес для шины Wishbone
 *   wb_we_o      - Сигнал записи/чтения (всегда '0' - чтение)
 *   pixel_data   - 8-битные данные пикселя, прочитанные из памяти
 *   data_valid   - Сигнал валидности данных на выходе pixel_data ('1' - данные актуальны)
 *
 * Протокол:
 *   При поступлении pixel_enable и если мастер свободен (не в цикле), мастер запускает
 *   транзакцию на шине (wb_cyc_o=1, wb_stb_o=1). Ждёт подтверждения wb_ack_i.
 *   При получении wb_ack_i завершает цикл и выдает данные на выход.
 */

module video_wb_master (
    input wire clk,
    input wire rst,

    // Интерфейс управления от видеоконтроллера
    input wire pixel_enable,
    input wire [23:0] phys_addr,

    // Wishbone Master Interface
    output reg wb_cyc_o,
    output reg wb_stb_o,
    output reg [23:0] wb_adr_o,
    output wire wb_we_o, // Постоянно '0', можно сделать assign
    input wire [7:0] wb_dat_i,
    input wire wb_ack_i,

    // Выход данных для видеоконтроллера
    output reg [7:0] pixel_data,
    output reg data_valid
);

    // Конечный автомат (можно реализовать и без явного FSM, как ниже)
    // Состояния: IDLE, REQUEST
    // Но в данном примере обойдемся регистром wb_cyc_o для простоты.

    // Логика работы
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            // Сброс всех выходных сигналов и состояний
            wb_cyc_o <= 1'b0;
            wb_stb_o <= 1'b0;
            wb_adr_o <= 24'b0;
            pixel_data <= 8'b0;
            data_valid <= 1'b0;
        end else begin
            // Снимаем строб по умолчанию (импульсный сигнал)
            wb_stb_o <= 1'b0;
            // Снимаем флаг валидности по умолчанию (импульсный сигнал)
            data_valid <= 1'b0;

            if (wb_ack_i) begin
                // Получено подтверждение от slave - транзакция завершена
                wb_cyc_o <= 1'b0;       // Завершаем цикл на шине
                pixel_data <= wb_dat_i;  // Защелкиваем пришедшие данные
                data_valid <= 1'b1;      // Сообщаем, что данные valid
            end
            // Если требуется пиксель и мы не находимся в середине транзакции...
            else if (pixel_enable && !wb_cyc_o) begin
                // Начинаем новую транзакцию на шине Wishbone
                wb_cyc_o <= 1'b1;       // Устанавливаем флаг цикла
                wb_stb_o <= 1'b1;       // Делаем импульс строба
                wb_adr_o <= phys_addr;  // Выставляем адрес на шину
            end
            // Дополнительная логика: если pixel_enable пропал во время транзакции,
            // мы все равно должны её завершить, дождавшись ack.
        end
    end

    // Мы всегда только читаем из памяти
    assign wb_we_o = 1'b0;

endmodule
