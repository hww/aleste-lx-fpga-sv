/**
 * Модуль: vid_addr_gen
 * Описание: Преобразует адрес CRTC (6845) в физический адрес видеопамяти.
 *            Поддерживает три режима адресации: Amstrad CPC, "Алеста" и линейный 32КБ.
 *            Добавляет базовый адрес из регистра для поддержки 24-битного адресного пространства.
 *
 * Входы:
 *   clk      - Тактовый сигнал (для возможной регистрации выхода)
 *   crtc_ma  - 14-битный адрес памяти от CRTC (Memory Address)
 *   crtc_ra  - 5-битный номер строки от CRTC (Row Address)
 *   mode     - 2-битный режим адресации:
 *                00: Режим Amstrad CPC
 *                01: Режим "Алеста" (чередование страниц)
 *                10: Линейный 32КБ режим
 *   page_reg - 8-битный регистр, задающий старшие биты адреса (базовая страница)
 *
 * Выходы:
 *   vram_addr - 24-битный физический адрес для видеопамяти
 *
 * Примечание: Реализация режима CPC является упрощенной и может требовать уточнения
 *             по документации на конкретный硬件.
 */

module vid_addr_gen (
    input wire clk,
    input wire [13:0] crtc_ma,
    input wire [4:0] crtc_ra,
    input wire [1:0] mode,
    input wire [7:0] page_reg,
    output reg [23:0] vram_addr
);

    // Внутренние сигналы для вычисленного адреса
    // Мы вычисляем младшие 16 бит, а старшие 8 берём из page_reg
    wire [15:0] internal_addr;

    // Комбинаторная логика преобразования адреса
    always @(*) begin
        case (mode)
            // Режим 00: Amstrad CPC (требует уточнения!)
            // В данном примере - простейшая реализация. Должна быть заменена на точную!
            2'b00: begin
                // !!! ВНИМАНИЕ: Это место требует перепроверки по документации на CPC!
                // Пример: старшие биты [16:14] формируются из RA[2:0], младшие - из MA.
                // Это предположение, а не точная реализация.
                internal_addr = { 2'b00, crtc_ra[2:0], crtc_ma[12:0] };
            end

            // Режим 01: "Алеста" (чередование страниц для четных/нечетных строк)
            2'b01: begin
                // Ключевой трюк: используем бит чётности строки (crtc_ra[0])
                // для переключения между верхней и нижней половиной 16КБ блока.
                // crtc_ra[0] = 0 -> Адрес в первой половине (0x0000 - 0x3FFF)
                // crtc_ra[0] = 1 -> Адрес во второй половине (0x4000 - 0x7FFF)
                internal_addr = { crtc_ra[0], 1'b0, crtc_ma }; // {A14, A13, MA[13:0]}
            end

            // Режим 10: Линейный 32КБ
            2'b10: begin
                // Простое линейное пространство: объединяем RA[0] и MA
                internal_addr = { crtc_ra[0], crtc_ma }; // {A14, MA[13:0]}
            end

            // default: на случай ошибки, используем режим "Алеста"
            default: begin
                internal_addr = { crtc_ra[0], 1'b0, crtc_ma };
            end
        endcase

        // Формируем окончательный 24-битный адрес:
        // Старший байт (A23-A16) из page_reg, младшие 2 байта - из internal_addr.
        // Выравниваем по границе 64K (page_reg * 65536) + internal_addr
        vram_addr = { page_reg, internal_addr };
    end

endmodule
